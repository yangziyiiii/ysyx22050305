module WBU(

);
    



    
endmodule //WBU

